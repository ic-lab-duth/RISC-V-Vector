localparam int SIM_VECTOR_INSTRS = 442;